netcdf run-mask {
dimensions:
	Y = 1 ;
	X = 1 ;
variables:
	int64 run(Y, X) ;
		run:_FillValue = NaN ;
	float lat(Y, X) ;
		lat:standard_name = "latitude" ;
		lat:units = "degree_north" ;
		lat:_FillValue = NaN ;
	float lon(Y, X) ;
		lon:standard_name = "longitude" ;
		lon:units = "degree_east" ;
		lon:_FillValue = NaN ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:source = "" ;
}
